<html>
<head>
<title>https://crecerjuntos.gob.sv/validate/certification/*H3T54P143130B5F79A5F7526437428G8S5D9C5F9</title>
</head>
<body bgcolor="#ebebeb">
<img src="images/verificacion.png" width="1340" height "600" align=middle">
